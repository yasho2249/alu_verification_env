program alu_tb();
   alu_env env ;
 initial 
       begin 
        env=new();
         env.run();
       end 
  endprogram        


